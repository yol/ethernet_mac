-- This file is part of the ethernet_mac project.
--
-- For the full copyright and license information, please read the
-- LICENSE.md file that was distributed with this source code.

-- Utility functions

library ieee;
use ieee.std_logic_1164.all;

package utility is
	-- Return the reverse of the given vector
	function reverse_vector(a : in std_ulogic_vector) return std_ulogic_vector;
	-- Extract a byte out of a vector
	function extract_byte(a : in std_ulogic_vector; byteno : in natural) return std_ulogic_vector;
end package;

package body utility is
	function reverse_vector(a : in std_ulogic_vector) return std_ulogic_vector is
		variable result : std_ulogic_vector(a'range);
		alias aa        : std_ulogic_vector(a'reverse_range) is a;
	begin
		for i in aa'range loop
			result(i) := aa(i);
		end loop;
		return result;
	end function;
	
	function extract_byte(a : in std_ulogic_vector; byteno : in natural) return std_ulogic_vector is
	begin
		return a((byteno + 1) * 8 - 1 downto byteno * 8);
	end function;
end package body;
